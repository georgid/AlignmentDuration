BZh91AY&SYx�6 & _�py���������`��� � �w� 2 z��a 4+"{`yBH6�A	@�I�xQ��j �44����d � ����� 2h� 2h�220CFi�F i�# ��RP�ѣI�10��F` )	�4�bjzM����=&jH�z�$��M!C�(i���= ����5�TVA�� @&
�
 U��^���W�4��v��)�@B�����\���H ��mɊ@ 8���>��#��OF���"��n]���湖=27N�� �J�^�nj��寱�ȥo��j�eQ2>�Pe�p�H� xx<{6li��Y�h-�zБ�4:�۲�YE�+�����wK�ڣJ��\hf���IWBSm����	n�@�D�3�7eK0�!����Vy�!<��y׫���I�L��%�%�N��ZJr�v�%�M����&m��v_N��0���f���-<�a����v�tN�����1�wΠ[l'{1��-�����^�{OOD�zO��}�d(�8��o1-knƦ͋pjlR�l�5u��mE��Lp�6RXl�a)T�5�-��a��[�Һ�H�a�K��mь�i-�X*"3R����-)GRl9ƱŐ��\�A�˴8Zյ�Ko�W^bԴ�"\G�W6��� �(�
 t��Һ�.�MMY���/��ⵜVqW�u������ʣjs�Sʦ8�$҄�Hς*�dɂ8H�!�L!��|��d�F�%��W���<��>�����/�x+j�[f�m�m,p9�\[�ˠ�K�WY73,�̻�M)ix�[[x�r�mSlF��R�BkV�).u
p��6�WH4��<�]-��v�\X]\ۈ�m�6s,�X���E\Ie��I�fn���`59c�M,
�,#vf��6k�6ز5�c�ƺ�8鯱�>���(���B+Q2=�Q��3X��h��@�	%S��"�U�����(+@��gE;S褜���?��o�D����F��%Y��v,!�Bq1�,)e�01�3г���t��ߕ�K��x��k�nf.����Z�*K���B���fbX��g�>¡Ӣ���-1d0���-
�M�֒��{�ӺDH�l @��oƆE����{` Z"j��0�%!$�%�����ݩF�1D�0��!��f�Y�-	:�Sot��zN��\���.�	iM309��)��q��.��2�����>񛪡��^s���0àd�b{�r����z�xf!���H��	mr&�UO�	��ID�o�1,6�����Q�C��w�v%�����ל���r�Wc�[�����..j���M�����]�)0���͈�s,� ����	퀐�$��5�"HN�x^��5&�	Z�I����������i"�LIw�S����k�s &�ff=���3b�+>=���gN�"�鼤���.yĄ8cg��� ���n�]H��%L.�q��*%0<�!�@�`�_�`��1C�rt�ZO�L�᳹��vF%C�Ï�؛�C���JٽR�`����<�y���ޛ������f<�'۔��ǌr���q�����֦)�<D���B ".��bCաl�T���{���[3s�zdʴ�%�|L{�D��cc�8���UV]r�+�+NR���S�H1b�\<�'�y���eu��j�w�;<=z��ژaF��vJ�2u	L�n��T�S:��;`�jնπ��(0n�}w���a.���6����������|�!�b|�Y|�Ja�z�ub$�gQ��q�31�ҞI���Վ�����}��"x=�(�g��]ϊ���^����O]B�ز{(�� �N�~�	��ދoɅ��0P�s�/o;9Z�mA-���~gW��%�RdZ�l���08�	���8F5�B�[o]�=w�z��z1�����`�h�-���3L��l6�<ɥ�!�,v��$�vg@ҙ��u:�z����o�t�|�=
�;~��Iy�|&{���q���S�i���ΆNE��r^���{���H&d���
JJeE�:��6���%��g��WT���=}�y�t�q�̹Q��o*^֟T�ӻ�zZ�o�u�rz�OHb�g�xK�DD�09Z�޼���򧢊N�޸%y\���_���m��SM�dQY9dt�oӎ0�j������{�ɥ��ʒ�G�=|��C{���׻���>� o�I|��b\wr"�C�-V:󐟀3���nݏ�����OS���^�[� �����\����4�G���GUf���J�%��%�M�K���ˉ�������3g��G [�y�{H���g�*~Tu�]�Rv`o2�:�U���A:�٭[�|�m�.>�f�G�DA�0�a����È�/��'����-����5��hԍ�4�RX����6&�k�ӒHNv���施��fff�m�n�� x^��塙�\��Z�Έ�'�g��	l�嘳f�W�/8)�f7�!$����`L������r��{�=��+�Kk�B�3���sj���.L2���]�c]�=��-��O�2���&dxJ'���R#�6,�M��v�mMEy�Y�]���0������t��U��үU)z�^�Ē�O�b��T�mxc��|Q�����;O��~U��p�	$�-4�PU RS���IO���w�%����tNr��-.��/��+��zV���f]�xn��X�3'�q���v�6�-_��o]븢����rSvj����yMt��E�L QPABRD�,'�:�fgRg$.K�	'pR��>�,�Gz1���!�L�pp�h�#��4�`�r��F]��98$^��c�5}������ķ�;�z>��O�^y>���9x��L����.9͝�����ˏ>F�҆�7�J	���q�q9�f"�k�a8��O��7-$�D
o��>�02�;bʆ�AP�1�|�����*��U�p�3% ���4�'=�e<��V�z��'<�wzc��s����^���{B/�*1aW�DXF<���	p@U`����s�3�ޞ�z�����Ҫ�H0�������%�L���7q�V����W��I0����L�e+;^\آ3�y�Mc0E�V�>��,gt݈���}�� �Un��b��:�5w��W���0�cAФ�%���)����a2]���_;�GO��_�5���_�c����.u&�a+����x�;��՜��= a�f���QUT���H�Ԃ�ϋ��%�@�O:�l*(*�����8� !*q��*Z�# B�J'�4#4����FNz�t��
J��Pj�һc��#���jpc��j�9�i ԻA�H�p*ClɁ�� �F"h&@�(����"JP�� �L��dh��JX��p�)
�v�ҩ%"L#��&�e!��K*T��G|켵�w�7q� �>D<�$B+"���H�g�e���W���mЙ_״A�2�D����}��u�	��w�R���n>�s�d/5��i���O
F�pϊtM�f��Q:/�2Xp?=��z,%	x�����Yy�W �6�q_�/���'�V��(+�	 D����(M134�Ad�𕨏̈́Cc���9}��C0�\I��٥O"�������݆_1%�O\2d�s �b��m������JfݍO�0k�}���q~r<�[�M&j]$ A @$�"D0����@ʤ�x 6�&"P�"��D��EkVa����5�3,2X^c^p�AQ��`f�D�Z��`�b=d^���x�����v���npw'�H����ux�C�+��LՄh|��w{��s?x��x��N6㭭� 0�T��o0`[��6=�_�6^�'�ߗU]�����+�d�He��r�}yI�1n.n>�:7;D�6���UU��}ϩ��F�J��9䐶G��-(��18�H"�XNa�p�!*� ��Thq�8� ��j�ZvAG��n�����ؐH�M�R�ȁ�-�
ѓ�Y��\)�j�
��X���p0U�
x���=��ˤ=�t�5N�I)Fu��n�a��uy��!A^��D#���w�

�wx�'�]�;�;�9T�AF! 4���l��pNc�;v|�����C��t,�-㴫[�2i(r���AA[Y���р�'�04$!,��`s��4} �0��#e�&#,�@YńL�L7��E~lyټÞ�D�¦"��Q�2�A�My&�9�>�>���.����Gs�4��
A��/�]��B@5��