BZh91AY&SY@,#X +�߀py���������`�e�  �v8�F�� � :��1 Bڀ��7�0@  � j$�H@ z��O)��@�4	*J4�4�2h2�	�@�4��d�L����L� ��IH( ���    �&��d�i�I�<���zC �h2)
h� �@    �gU@BA��PT&��7 ��v�����AB�'�;����CJ�a'��UX��B�����Z�D
����d�pv���[ݻ�� ������F�[��*rZ)OS+�K�b_
ʼi�rNnm�v<�������N��,����(�럾��p���i��������K�{�;�<�����ѷeԲ�lW��<�'9���'ux���mQ�Jnܺ�(uÒUД�A'�M��<8Kv��
&�9�(�a Cq{;x���]�p�<�������L��%�%�N��ZJr�v�%�M����&m��v_N��0���f���-<�a����v�tN�����1�wΠ[l'{1��-�����^�z���C�{��x���
;�jq�����cSfŸ56)ev�Ӻ=u��ZK��X�;;��ݺ]�M�:�s�v��N��܅�G���]�Uc{3ڝH�u�	��^�ۮ�����\��*�Q�w3B��:٩��ٝ���qgH2��7C��e�����])�ײ�;��u��z�U�f�����z���lj��]�	f@�b{���d:uc7T-�}�/�Eq�x������d���h�8Ъ�΂�k�"�$�X0�15����~p�(#��үC�S)D�H fD#�0Hd�dS)`zN�b'�ۚ[�n��3}B�r�((6�0�2SnSi`ˁ�r���]�]
�ɹ�f�e�jiKK�����ś��j�b5�P��JZ��Is�S�i���A�/��͚�o &K�"�����F�mI�Ø!frĄXm�*�K-��M[3t�g����i`W9a��41�V͠�����[K��2��m�t���A�J�/= ��~��B�h�"��	%R���"U������	0�|2����'4Ԙ�B' Hٿ��At�.�I�Y�<*�'�'#"^#�*&D
��N#�1/vd�*U��b�M#\��0�'&���:�1$�,H��ۙ��s���Ɩ�
��B0ĸ�X q`��!lk̺Bڙ4D�18���ݿ/���dQ��~>�'��)l���4D�@ ���w�4*�%i��f�Y$3������2B�{,��3��
s �z 1 C��׺�{n�ũD��ގ�sC}V3��
�.�%q���T�(�6���r�k�2f�.�; @]�7OPx�i83���ب�A�o��Qv�љ�"A!ڍpl�)iɀ ;��y��d;�j�y� zX���ݻ�V��k3Y�E�e�2%E�Ҁ�$[��@� zw�0���kS}�@��>�s��7-��}��" `��jр F�����3�n��N�H}����32�$�!H��ǌQ��eyT����.fb  �*���޸On�U������Xs�"� dD@�a��0�����(?������C��	�D焖�E�8���b,�ٽ��^������ƺ��J�]�kX��İu�I?�� ~6�L�����t좑f�R�a����6��	3+?��.��d/{;��G��ߠ�Y��T)琰���Њ�H��ɮȈ xUnQ�3�7>����� �#]��L��
h̐ d��$�U�qTg��g~a x��"pkc*�D��|@��%��ź�p�*n2�����Wy�\�+�q�$1�(�Nd0S��2���l��oR��4��)W���4� �8ǡՠ̌Ǥ�9&� x�@�S]u�[c���6�ӰC� n� v<���KMH���0	�b rcż9�	�r廝� W*f~l#(K4V^RŜ�с�ª_!�����>�D@���Яz�F�J:�Ժ8F�e,d{��'=���X]x��A%��L�,xڧ�O���+k�����C������H�\ 
��JǔP��_z�|�� �Vdg� �����u|�8TzJ1p��}z�;X�" p$,)B@2Й������\�`�h/-�qv�.�9�k����%0���n24X��H�������$�a ��\~��3sa��k��3V-����7�7oM���i�z|A4��"�6r���o@�/*�7�^�^�ɪa62�H�Z�<ę2�-��ںz�Z��c^(��h#F��5n@���f�m�p؈<h� ��<lt?S�)(O���Z����L��5GƀҸ:0�T�̄Dˣ0 &D����׎L�R��R�����b����_:cpY�0e"$�Q"�$	¬ֶ��k!��`� ���;��'���Y�BA_�TG�c�׻��q{��V�ߔ g�J��b|�r�IWʪ�q��٭G�'��� ml�F"�.���	*���  /m���D�u��O�	�=�����N�{#��V�&��i�-"�3��+���7j����|s�c�þ=> 	�yo��Wz�M?�z�����Q E���7�ܞ�F���vg��� Q���H��" ĉN0���RDa�Q��z�잞x�4k�[	Aa�kI�ѩ2(i������lL�.X$�Q��@ !ゎ���~�&eZ3Q�.���L�[����I���Q䄑�C��M�o=<^���{��g��Ú��ލ�qe);�D X��'�L)SH�0k����0���g/�k�W���d�z&+ޗ���3��p$�1�o��~yc� �z R�\�  ���?T�3�3-��T�mXb�F{���F��v�U���4noˍP�O  EO��u��U�Iy���^��Su'�64�kFZ�$� �m������ʔTFj�g��/5��S3�y��I�A�&	�R����$ ��8κ��>h��U�ld��2G���^�̲O�ύ.s� ܺ��oёOq#���]�~�a��z^#��׻rcCN͚�ޱ���B�a��j��s�64��u�L��\�.7�9$TP��5�	�}�,�����fm�,�yH�A	���Q56V{�t����,-;pp�h�#��4�`�r�,!,��0�,��&�=�P�-�R�A2�A�s���/{��F��(��mIK<~Lx� #V&ñ��h��*py�7�N'�=D$s9׳�k��DC"4���2	\0�
B{0�����C�uemߣ���E*�&C�� �\;u�\8���J�/0@��U���T�3N�r�[��8��&��A-I� �T˿�����3<u�O|r�]Ѫ���#����"@�%	R�R�X@U��"� BAX �0x� ���'�WxJۥ7��n���=<�uy�n4I�'}�~�8��og����� 	&'�;P�#UTyf��oV��.��#�#�� 	���B����z]Yyz)��7� @��O��Ӫ�n���W{�4�"(�b &�%�	2�M@ee��с�v&_~s���o]�|��Nh���2滦�j���E������DDR�O���̷���@~S��D��TQT���� � 8r'JyA�5�
h�*>�LN8�f
'�0`[֭ EslV*D S
@�����3KJ�# ,��%�(Y^�Md�DBJ˒ `0�j5�@�ˠ���R�RG��	S+E�'h6(�PL<o7��%��l�9�Fj�I5Rsf�ެu&��o,L'l�!�FK`I�e�JFF&T�	�!��4��I(Fa)V�A�Ѭ�2"6��,��Gl�z�8� ����^�(A)J!��|)t�R1�e�<�����Od��bj��`:P?*{�����2�g�e���y�0�g��^u�6a��Jl��t2Oe�!�`K����}�9FD������,��@�^F����C� ���4�U��D�zG�ú(M5�R�H0�$��ej#�$��g�ìy�vx*����G�a�-� �5��6F��h�����a$�O:iU��JU��U�����ga����I��+�?��ӓ��G~})t��t���A �$��(2C
H� J�w�C 7�L(��2"��E�EkT��J%��VJB���G�(��l(MA����ۛ�'i9�D�Ѳ2Z�j���w�;�H;=��u4��� 0M���L[x����\���]�Z���cP�y4��yN�,}e�����u�<���j��T.HC(Q��Iq�ve����qr\}p�� �����Gz����>�H��S�zd��C�4KJ(�MN�t����TO7SA��C�� 
�8���7��6<�9ɺ�ZQM����&
<)�<�)#x�I�V�� NH�J��I:v�������Ȫ�o�,Q�����"�����>&���?T�P3Q��J1\�7�m1$�y�6��T�`�+����_�U����.ۊi0�*�B��dX�Ay���P�@M�X��;��t��ay`���'9T��ՙ5�%�~~QЪ�Z�u��8-�&���aYc!�fgN�����df�-�0�BW���!G�B`��H?�;��cM@�HQ�UP<Jؚ�Ih !�5�5��
a?pYl�hj�Aؒ�4N#�H�K�w$S�	�5�