BZh91AY&SYS��� 1v_�ppy���������`�|��  �ܠ�9.��4� 4�  � ^��  4@H�d4  �ѓMi� ��$�%=M4�4��26�  dɣ��i�0LM4����RDR����z� 14�  "QA&&����@�~�ɦ��O(������P�M     ��T)ȣҠ�DUΪ�m�|��7�����0�)Q��s��AE�DA#	�UUUW$
��B��I��%�TK���;�/o�P��Y�o����� �-�Xu���/ʅ/����`[G�om�����UiuS0c������bg �E+4ȑ�A�}P�\���:��?��_� �N��7���C�>�s�M�O_O����76�BM\Kv�V���I���p�z8py�^���^.�2�5ݺ�Z���%�	]�����n��ݸ�)��1�4�7J�S1w$���!���)���ɤ�}��tO(_ٻX�3�*W�۵��^X�n�e�Dʛu�����A�d�q��l8�����0�[Y�t�{8n����O=y��<��֪�[lR׃{a���??>c���/�����y�ί%��l�ݝ]�$�uvkJ���^�wY{3�\�9�at�Ԝ���\0�F�{	Xi�Y7n����u��Ft��57a�$!zi�ĝ�vPc��Xv�ۮ:R�.�;54��[ ��D�s�#�ޕ;)��!�^�C�gg]I�tD�kG���NaS#;){�㬳M��-�A��B�s�&����wQ!�N����;�D�s�e%$�N������H]Ժ�+�MMY���-I,�$�	�'9:Qs�;�~Jd�Q.a���-� ]"8k�M��s0GF��R��1�8��h�G�~r��u�K�I��ل�֪		AF!JB�s��H!�A0�D0���秝�'�{V��B\���|빹ׅ�_��ez�I�i��ܮ�\�K4��MˆL��j��4������]���HnWX�XR��B����E.��x��6Գ+��L�0�Y�x�hݪI�7Y��%�ڦ�ei�"$��I3�R��YM.54����b�f�A!m2��SaRʩh$E��)Y���@��V)��@g�LU И��K���Zd^P�a�s������[D #`	GDU"/�5����R� ���d��p��C�e�T)�V���v[��⟬Nӗ�d��;�kz�٢9�NF$'# ֗��α4�Ӈ^m�K0�|u֚@�Y��Q-D!���4�Iń�`��� E��W�4�;�z�պGM"��ͷC7]&�f��ų��%<���jff��� �7ĜYe8�r���IR rwRAC�J		%+J9j���->������Jr�c��mN�H���$Skl~��������#����:��4��V��}�fJ���˟��o�w�:w^4s�`i:�s�vJ��7	Ƭd�:[L��x�N�&(�'��:���N9w��	G
Z��r�%:S&���IW�y�d���vh���P�U���]8�����
�㳮hym�(f�
A��m�8�E�?+��},��;_%׮Q7B��:e0z%��m�ۺ�}.�����*�p�p�.��Ġ�T#	Ǒ3��=�i	�^�_^g���ܕ蕜�[�����x�n!����]�)0�{��ۙ��7�&�0��'�B�(��4��"HN�x^���f�%i�=Bw�������!���{������&�J���xu�c6v��a�(� ]��ǻ]�`a�YwO�����x]ìq��f`�G(�����Nr"<Z����}��K'\�w%��[�ɈL�E͊�L��4f�+�����y����S��<�w�dk՗yCsk�v��sin��0ҡ���m6�sh{;�[7�̹<��Mfס�*s�X-vf�&�
�A�1���ȣ���&<UnR�31ʋ�Uƴ8��p�6mDS�x�˨��̈�]5�����ٚ�Gaa�����0
i�ӽ���t,6d�-3����a���7]���p�9����%�,{a���L�aԜ�a�ۿ�s�zy�y덏�5��0������_A �]٘4L�g��{�ژi+$�IV�3'P��~Jq���2R)�5�Kjg3����è�D@Ѹ�0�z�!��P�v���]��3D68�-������mT�J�������"U'��~T����yj&־.E�eǨ�31�%QW�h�5c�s7��&��HA���-D��B �tz�����+�ݡ�I��&�F=OmI��~@0մ}>4.ݸ&�v�ACϺa6�Q��=�p���W_z��ϫ��D/��º��u|����Q<__���ȶ�f&Ԃ �#₤�	aA��ϭO��)���s�x���[k3v�n14�[1���Ѯc��ې��/*<�����:`^��p��$�����C�D�����>�<�>�w:���3c���A��0�'g�.ç�4���*ʺѮ`�*�m�3m��)��mɄ��`� �TGI
�S*0�u8J�vX�%��xԨuJ�K�����"�s1\k3.T#X�
E��l��>��jwu>�kAo�0��qqT�P��k^)Zi�xJT��v	���}y�ȃ秂�d�w�J^e�W�׻kff�5-lJ)	2L������:�k�y�,N$Bmu:���������微��vY�q�'�Sצa�u�f��䮭?& �/Oyǘ���L���?�j���A<Q^f����NM�?��DÐ-zz��|� ar�K��]��o��=�{Z�˸LN�jW�7�f�u8�
��E("^]�]���T��wm�#M���������f!�����'�>��Qow��?Tu����'�^)36od.N��W˹�Y�K[}�L�� ���,"D�qcXI�0�F##�~!�;�	�e�6�VAؖT�ı%4d\jT��;M�)��E��!�� 1˦LK|9��vOSOp�����Rӯ
	���C���{�F�y܄36s�����\磍g	�����Zq�0�lҊ�͹�>���me��BIu�3�Ď(-뼿i�(���Ȉ̳޷��H�6�t�r�;@W�D�}]#��h�2�&�x<�T��Ճ>C�;��	�lG"}Q�2 �U
"fY�¡T��!]���V6'4�ٱC�n�z���G�����ʯ+|�Egdf��'=��K�ki4��^���kjIV�o�V!*)�U*dm��xB��∈xt�k���v{'��/��sZ�3���I�M%P�I�&
X`$��a�DaE`�́k*n���������Gg�O��+��g�o2y���;�<�ZP��W�V*���+�����!���6���z�̾ �^Jc�mX�wn��(�S�ks�e��H(� �)"��-��|�B�I>��	�����(�Q&��
"b�y��|�'��ᮚܼY�Y"2�8���f����Wzx$L2�X�I�xD�>�}�TƉ*���_3�=�>eK�!�QN��(�+xMII-���;��`�$��ҩ2�i�KAqg�ڐ���H�C���>ܟ��3GC4���l�(!KI.���s�f"�k҇�|W����w�E�J�D=g%�a��qۤ�XKx�$�v�f}0;�����H�y�T���I��we �8�&��/�8��^�6��ϮG�-�H��l�T��,��U��a���=�����NH������,��e�abf8ID�TM�ff8�'�vq8�fN[��sw+ſ����oS娨��.�x�O�r]$��1|7q�V�˜�>� $�	#��5SL���\Fh�M&ts��x�$qN�k�-�[�S�Q<�S�4Z��T���=�l�A��5��֓<�����m��֙�L����\xRH��wyviO������v�D��}���;4��;��f��W�;e�wFq��йԛvN�	�9���b�^<{lW|�����yf�i�ꪦ���$D�R�!ӱz�[���q}�m� ��ј*��0bY ��0��P�a�R(�!��J�1#,��� �E+�S��	/=���VÌ�s�@�4m�"�8 j� =x�o8!��3�C�W�Wfj^<uo8k��Vs�ÆueNN��/���a1�.�fPaa�!�b`R��D,IA�8H�P�H�R��B�H�-)� �()ZEݕ�J�%*�*n@a�HkXDl��p��&"��&���	e!?�`z(v�@�Ȉ�Q$D��Pe�G�O)��av����O�P�n]m��"*X!<��6<���Q����6W!��k����=�v�g:�ܻ���~�f���m�#������%�AuA���[��ן/���l��Q5I$��-�b�fkѸ����'ҁ���	�<�DD�aO�f�	aT�h=���+EO8��#Q���j�E��DA.���ϟ�E�=�\��U�_UZo���$���x@#���-��
�,���PN9m�X�Ma�-�I B����ӂ��a�2Y�)��"b����A �$�C �2�$2��,'z�R af
��`"��D7n8ܲ�౸8١`��0��J�!����*mn��Ɉl��\�Pbf�1��*�O����iq؇x1����~����0QԻ��!Pym ;9ð���� �Nt�i�on��V�à��C!�[_����7�o���?%ýӀ�q��4REh-;?��'㜯q�p0�<�0�^i ��AE�y�Oc�����/.N��b����Ŋ��@�@���o��D� ���K��TN��9�������\�r�j�ZD`�T~��� �BպoHP��`�.B�]��nDA,:9NY��9z���'?ij��ҹ*��'����~�y��/���Z���Rj\}��ň'qD�<�^QN��Y:����Z��Z}�=j]K�;�H��h����E�R<��"PC0���-Xn=<}�8s��ɟH���u�5*�"���^Ä�^�� i�"�4"�\�P���P���c��E
���j_B�j�3�J��0FE���] k��D��Ư uY�\�v  �h]j��&EWu@��A>Vi�~F��`�Ц��J�A� �=8���rE8P�S���